magic
tech gf180mcuD
magscale 1 10
timestamp 1757535624
<< nwell >>
rect -2080 60 -800 452
rect -2080 -120 -740 60
<< pwell >>
rect -20 -920 2356 -640
rect 2480 -920 4856 -640
rect -13480 -2200 -9984 -1920
rect -6580 -31940 -5908 -3224
rect -5780 -31940 -5108 -3224
rect -4980 -31940 -4308 -3224
rect -4180 -31940 -3508 -3224
rect -2580 -31940 -1908 -3224
rect -1780 -31940 -1108 -3224
rect 1220 -31940 1892 -3224
rect 2020 -31940 2692 -3224
rect 2820 -31940 3492 -3224
rect 3620 -31940 4292 -3224
rect 5220 -31940 5892 -3224
rect -6380 -33000 -6100 -32080
rect -5580 -33000 -5300 -32080
rect -4780 -33000 -4500 -32080
rect -2380 -33820 -2100 -32076
rect 1420 -32760 1700 -32064
rect 2220 -32760 2500 -32064
rect 3020 -32760 3300 -32064
rect 3820 -32760 4100 -32064
rect -6580 -62640 -5908 -33924
rect -5780 -62640 -5108 -33924
rect -4980 -62640 -4308 -33924
rect -4180 -62640 -3508 -33924
rect -2580 -62640 -1908 -33924
rect -1780 -62640 -1108 -33924
rect 420 -62600 1092 -33884
rect 1220 -62600 1892 -33884
rect 2020 -62600 2692 -33884
rect 2820 -62600 3492 -33884
rect 3620 -62600 4292 -33884
rect 5220 -62600 5892 -33884
<< nmos >>
rect 48 -808 2288 -752
rect 2548 -808 4788 -752
rect -13412 -2088 -10052 -2032
rect -6268 -32932 -6212 -32148
rect -5468 -32932 -5412 -32148
rect -4668 -32932 -4612 -32148
rect -2268 -33712 -2212 -32144
rect 1532 -32692 1588 -32132
rect 2332 -32692 2388 -32132
rect 3132 -32692 3188 -32132
rect 3932 -32692 3988 -32132
<< ndiff >>
rect 48 -677 2288 -664
rect 48 -723 61 -677
rect 2275 -723 2288 -677
rect 48 -752 2288 -723
rect 2548 -677 4788 -664
rect 2548 -723 2561 -677
rect 4775 -723 4788 -677
rect 2548 -752 4788 -723
rect 48 -837 2288 -808
rect 48 -883 61 -837
rect 2275 -883 2288 -837
rect 48 -896 2288 -883
rect 2548 -837 4788 -808
rect 2548 -883 2561 -837
rect 4775 -883 4788 -837
rect 2548 -896 4788 -883
rect -13412 -1957 -10052 -1944
rect -13412 -2003 -13399 -1957
rect -10065 -2003 -10052 -1957
rect -13412 -2032 -10052 -2003
rect -13412 -2117 -10052 -2088
rect -13412 -2163 -13399 -2117
rect -10065 -2163 -10052 -2117
rect -13412 -2176 -10052 -2163
rect -6356 -32161 -6268 -32148
rect -6356 -32919 -6343 -32161
rect -6297 -32919 -6268 -32161
rect -6356 -32932 -6268 -32919
rect -6212 -32161 -6124 -32148
rect -6212 -32919 -6183 -32161
rect -6137 -32919 -6124 -32161
rect -6212 -32932 -6124 -32919
rect -5556 -32161 -5468 -32148
rect -5556 -32919 -5543 -32161
rect -5497 -32919 -5468 -32161
rect -5556 -32932 -5468 -32919
rect -5412 -32161 -5324 -32148
rect -5412 -32919 -5383 -32161
rect -5337 -32919 -5324 -32161
rect -5412 -32932 -5324 -32919
rect -4756 -32161 -4668 -32148
rect -4756 -32919 -4743 -32161
rect -4697 -32919 -4668 -32161
rect -4756 -32932 -4668 -32919
rect -4612 -32161 -4524 -32148
rect -4612 -32919 -4583 -32161
rect -4537 -32919 -4524 -32161
rect -4612 -32932 -4524 -32919
rect -2356 -32157 -2268 -32144
rect -2356 -33699 -2343 -32157
rect -2297 -33699 -2268 -32157
rect -2356 -33712 -2268 -33699
rect -2212 -32157 -2124 -32144
rect -2212 -33699 -2183 -32157
rect -2137 -33699 -2124 -32157
rect 1444 -32145 1532 -32132
rect 1444 -32679 1457 -32145
rect 1503 -32679 1532 -32145
rect 1444 -32692 1532 -32679
rect 1588 -32145 1676 -32132
rect 1588 -32679 1617 -32145
rect 1663 -32679 1676 -32145
rect 1588 -32692 1676 -32679
rect 2244 -32145 2332 -32132
rect 2244 -32679 2257 -32145
rect 2303 -32679 2332 -32145
rect 2244 -32692 2332 -32679
rect 2388 -32145 2476 -32132
rect 2388 -32679 2417 -32145
rect 2463 -32679 2476 -32145
rect 2388 -32692 2476 -32679
rect 3044 -32145 3132 -32132
rect 3044 -32679 3057 -32145
rect 3103 -32679 3132 -32145
rect 3044 -32692 3132 -32679
rect 3188 -32145 3276 -32132
rect 3188 -32679 3217 -32145
rect 3263 -32679 3276 -32145
rect 3188 -32692 3276 -32679
rect 3844 -32145 3932 -32132
rect 3844 -32679 3857 -32145
rect 3903 -32679 3932 -32145
rect 3844 -32692 3932 -32679
rect 3988 -32145 4076 -32132
rect 3988 -32679 4017 -32145
rect 4063 -32679 4076 -32145
rect 3988 -32692 4076 -32679
rect -2212 -33712 -2124 -33699
<< pdiff >>
rect -1894 253 -1768 266
rect -1894 79 -1881 253
rect -1835 79 -1768 253
rect -1894 66 -1768 79
rect -848 66 -800 266
<< ndiffc >>
rect 61 -723 2275 -677
rect 2561 -723 4775 -677
rect 61 -883 2275 -837
rect 2561 -883 4775 -837
rect -13399 -2003 -10065 -1957
rect -13399 -2163 -10065 -2117
rect -6343 -32919 -6297 -32161
rect -6183 -32919 -6137 -32161
rect -5543 -32919 -5497 -32161
rect -5383 -32919 -5337 -32161
rect -4743 -32919 -4697 -32161
rect -4583 -32919 -4537 -32161
rect -2343 -33699 -2297 -32157
rect -2183 -33699 -2137 -32157
rect 1457 -32679 1503 -32145
rect 1617 -32679 1663 -32145
rect 2257 -32679 2303 -32145
rect 2417 -32679 2463 -32145
rect 3057 -32679 3103 -32145
rect 3217 -32679 3263 -32145
rect 3857 -32679 3903 -32145
rect 4017 -32679 4063 -32145
<< pdiffc >>
rect -1881 79 -1835 253
<< psubdiff >>
rect -6556 -3320 -5932 -3248
rect -6556 -31844 -6484 -3320
rect -6004 -31844 -5932 -3320
rect -6556 -31916 -5932 -31844
rect -5756 -3320 -5132 -3248
rect -5756 -31844 -5684 -3320
rect -5204 -31844 -5132 -3320
rect -5756 -31916 -5132 -31844
rect -4956 -3320 -4332 -3248
rect -4956 -31844 -4884 -3320
rect -4404 -31844 -4332 -3320
rect -4956 -31916 -4332 -31844
rect -4156 -3320 -3532 -3248
rect -4156 -31844 -4084 -3320
rect -3604 -31844 -3532 -3320
rect -4156 -31916 -3532 -31844
rect -2556 -3320 -1932 -3248
rect -2556 -31844 -2484 -3320
rect -2004 -31844 -1932 -3320
rect -2556 -31916 -1932 -31844
rect -1756 -3320 -1132 -3248
rect -1756 -31844 -1684 -3320
rect -1204 -31844 -1132 -3320
rect -1756 -31916 -1132 -31844
rect 1244 -3320 1868 -3248
rect 1244 -31844 1316 -3320
rect 1796 -31844 1868 -3320
rect 1244 -31916 1868 -31844
rect 2044 -3320 2668 -3248
rect 2044 -31844 2116 -3320
rect 2596 -31844 2668 -3320
rect 2044 -31916 2668 -31844
rect 2844 -3320 3468 -3248
rect 2844 -31844 2916 -3320
rect 3396 -31844 3468 -3320
rect 2844 -31916 3468 -31844
rect 3644 -3320 4268 -3248
rect 3644 -31844 3716 -3320
rect 4196 -31844 4268 -3320
rect 3644 -31916 4268 -31844
rect 5244 -3320 5868 -3248
rect 5244 -31844 5316 -3320
rect 5796 -31844 5868 -3320
rect 5244 -31916 5868 -31844
rect -6556 -34020 -5932 -33948
rect -6556 -62544 -6484 -34020
rect -6004 -62544 -5932 -34020
rect -6556 -62616 -5932 -62544
rect -5756 -34020 -5132 -33948
rect -5756 -62544 -5684 -34020
rect -5204 -62544 -5132 -34020
rect -5756 -62616 -5132 -62544
rect -4956 -34020 -4332 -33948
rect -4956 -62544 -4884 -34020
rect -4404 -62544 -4332 -34020
rect -4956 -62616 -4332 -62544
rect -4156 -34020 -3532 -33948
rect -4156 -62544 -4084 -34020
rect -3604 -62544 -3532 -34020
rect -4156 -62616 -3532 -62544
rect -2556 -34020 -1932 -33948
rect -2556 -62544 -2484 -34020
rect -2004 -62544 -1932 -34020
rect -2556 -62616 -1932 -62544
rect -1756 -34020 -1132 -33948
rect -1756 -62544 -1684 -34020
rect -1204 -62544 -1132 -34020
rect -1756 -62616 -1132 -62544
rect 444 -33980 1068 -33908
rect 444 -62504 516 -33980
rect 996 -62504 1068 -33980
rect 444 -62576 1068 -62504
rect 1244 -33980 1868 -33908
rect 1244 -62504 1316 -33980
rect 1796 -62504 1868 -33980
rect 1244 -62576 1868 -62504
rect 2044 -33980 2668 -33908
rect 2044 -62504 2116 -33980
rect 2596 -62504 2668 -33980
rect 2044 -62576 2668 -62504
rect 2844 -33980 3468 -33908
rect 2844 -62504 2916 -33980
rect 3396 -62504 3468 -33980
rect 2844 -62576 3468 -62504
rect 3644 -33980 4268 -33908
rect 3644 -62504 3716 -33980
rect 4196 -62504 4268 -33980
rect 3644 -62576 4268 -62504
rect 5244 -33980 5868 -33908
rect 5244 -62504 5316 -33980
rect 5796 -62504 5868 -33980
rect 5244 -62576 5868 -62504
<< nsubdiff >>
rect -2056 356 -800 428
rect -2056 -24 -1984 356
rect -2056 -96 -740 -24
<< polysilicon >>
rect -5600 -740 -5480 -720
rect -5600 -820 -5580 -740
rect -5500 -760 -5480 -740
rect -540 -740 -420 -720
rect -540 -760 -520 -740
rect -5500 -800 -5400 -760
rect -600 -800 -520 -760
rect -5500 -820 -5480 -800
rect -5600 -840 -5480 -820
rect -540 -820 -520 -800
rect -440 -820 -420 -740
rect -540 -840 -420 -820
rect -180 -740 -60 -720
rect -180 -820 -160 -740
rect -80 -760 -60 -740
rect 4880 -740 5000 -720
rect 4 -760 48 -752
rect -80 -800 48 -760
rect -80 -820 -60 -800
rect 4 -808 48 -800
rect 2288 -808 2332 -752
rect 2504 -808 2548 -752
rect 4788 -760 4832 -752
rect 4880 -760 4900 -740
rect 4788 -800 4900 -760
rect 4788 -808 4832 -800
rect -180 -840 -60 -820
rect 4880 -820 4900 -800
rect 4980 -820 5000 -740
rect 4880 -840 5000 -820
rect -5600 -1180 -5480 -1160
rect -5600 -1260 -5580 -1180
rect -5500 -1200 -5480 -1180
rect 4896 -1180 5016 -1160
rect 4896 -1200 4916 -1180
rect -5500 -1240 -5400 -1200
rect 4800 -1240 4916 -1200
rect -5500 -1260 -5480 -1240
rect -5600 -1280 -5480 -1260
rect 4896 -1260 4916 -1240
rect 4996 -1260 5016 -1180
rect 4896 -1280 5016 -1260
rect -9960 -2000 -9860 -1980
rect -13456 -2088 -13412 -2032
rect -10052 -2040 -10008 -2032
rect -9960 -2040 -9940 -2000
rect -10052 -2060 -9940 -2040
rect -9880 -2060 -9860 -2000
rect -10052 -2080 -9860 -2060
rect -9620 -2000 -9520 -1980
rect -9620 -2060 -9600 -2000
rect -9540 -2040 -9520 -2000
rect -9540 -2060 -9420 -2040
rect -9620 -2080 -9420 -2060
rect -10052 -2088 -10008 -2080
rect 6220 -2740 6260 -2640
rect 6160 -2760 6260 -2740
rect 6160 -2820 6180 -2760
rect 6240 -2820 6260 -2760
rect 6160 -2840 6260 -2820
rect 6160 -2920 6260 -2900
rect 6160 -2980 6180 -2920
rect 6240 -2980 6260 -2920
rect 6160 -3000 6260 -2980
rect 6220 -3060 6260 -3000
rect -6344 -3473 -6144 -3460
rect -6344 -3519 -6331 -3473
rect -6157 -3519 -6144 -3473
rect -6344 -3582 -6144 -3519
rect -6344 -31645 -6144 -31582
rect -6344 -31691 -6331 -31645
rect -6157 -31691 -6144 -31645
rect -6344 -31704 -6144 -31691
rect -5544 -3473 -5344 -3460
rect -5544 -3519 -5531 -3473
rect -5357 -3519 -5344 -3473
rect -5544 -3582 -5344 -3519
rect -5544 -31645 -5344 -31582
rect -5544 -31691 -5531 -31645
rect -5357 -31691 -5344 -31645
rect -5544 -31704 -5344 -31691
rect -4744 -3473 -4544 -3460
rect -4744 -3519 -4731 -3473
rect -4557 -3519 -4544 -3473
rect -4744 -3582 -4544 -3519
rect -4744 -31645 -4544 -31582
rect -4744 -31691 -4731 -31645
rect -4557 -31691 -4544 -31645
rect -4744 -31704 -4544 -31691
rect -3944 -3473 -3744 -3460
rect -3944 -3519 -3931 -3473
rect -3757 -3519 -3744 -3473
rect -3944 -3582 -3744 -3519
rect -3944 -31645 -3744 -31582
rect -3944 -31691 -3931 -31645
rect -3757 -31691 -3744 -31645
rect -3944 -31704 -3744 -31691
rect -2344 -3473 -2144 -3460
rect -2344 -3519 -2331 -3473
rect -2157 -3519 -2144 -3473
rect -2344 -3582 -2144 -3519
rect -2344 -31645 -2144 -31582
rect -2344 -31691 -2331 -31645
rect -2157 -31691 -2144 -31645
rect -2344 -31704 -2144 -31691
rect -1544 -3473 -1344 -3460
rect -1544 -3519 -1531 -3473
rect -1357 -3519 -1344 -3473
rect -1544 -3582 -1344 -3519
rect -1544 -31645 -1344 -31582
rect -1544 -31691 -1531 -31645
rect -1357 -31691 -1344 -31645
rect -1544 -31704 -1344 -31691
rect 1456 -3473 1656 -3460
rect 1456 -3519 1469 -3473
rect 1643 -3519 1656 -3473
rect 1456 -3582 1656 -3519
rect 1456 -31645 1656 -31582
rect 1456 -31691 1469 -31645
rect 1643 -31691 1656 -31645
rect 1456 -31704 1656 -31691
rect 2256 -3473 2456 -3460
rect 2256 -3519 2269 -3473
rect 2443 -3519 2456 -3473
rect 2256 -3582 2456 -3519
rect 2256 -31645 2456 -31582
rect 2256 -31691 2269 -31645
rect 2443 -31691 2456 -31645
rect 2256 -31704 2456 -31691
rect 3056 -3473 3256 -3460
rect 3056 -3519 3069 -3473
rect 3243 -3519 3256 -3473
rect 3056 -3582 3256 -3519
rect 3056 -31645 3256 -31582
rect 3056 -31691 3069 -31645
rect 3243 -31691 3256 -31645
rect 3056 -31704 3256 -31691
rect 3856 -3473 4056 -3460
rect 3856 -3519 3869 -3473
rect 4043 -3519 4056 -3473
rect 3856 -3582 4056 -3519
rect 3856 -31645 4056 -31582
rect 3856 -31691 3869 -31645
rect 4043 -31691 4056 -31645
rect 3856 -31704 4056 -31691
rect 5456 -3473 5656 -3460
rect 5456 -3519 5469 -3473
rect 5643 -3519 5656 -3473
rect 5456 -3582 5656 -3519
rect 5456 -31645 5656 -31582
rect 5456 -31691 5469 -31645
rect 5643 -31691 5656 -31645
rect 5456 -31704 5656 -31691
rect -6260 -31960 -6160 -31940
rect -6260 -32020 -6240 -31960
rect -6180 -32020 -6160 -31960
rect -6260 -32040 -6160 -32020
rect -5460 -31960 -5360 -31940
rect -5460 -32020 -5440 -31960
rect -5380 -32020 -5360 -31960
rect -5460 -32040 -5360 -32020
rect -4660 -31960 -4560 -31940
rect -4660 -32020 -4640 -31960
rect -4580 -32020 -4560 -31960
rect -4660 -32040 -4560 -32020
rect -3860 -31960 -3760 -31940
rect -3860 -32020 -3840 -31960
rect -3780 -32020 -3760 -31960
rect -3860 -32040 -3760 -32020
rect -2260 -31960 -2160 -31940
rect -2260 -32020 -2240 -31960
rect -2180 -32020 -2160 -31960
rect -2260 -32040 -2160 -32020
rect -1460 -31960 -1360 -31940
rect -1460 -32020 -1440 -31960
rect -1380 -32020 -1360 -31960
rect -1460 -32040 -1360 -32020
rect 680 -31960 780 -31940
rect 680 -32020 700 -31960
rect 760 -32020 780 -31960
rect 680 -32040 780 -32020
rect 1480 -31960 1580 -31940
rect 1480 -32020 1500 -31960
rect 1560 -32020 1580 -31960
rect 1480 -32040 1580 -32020
rect 2280 -31960 2380 -31940
rect 2280 -32020 2300 -31960
rect 2360 -32020 2380 -31960
rect 2280 -32040 2380 -32020
rect 3080 -31960 3180 -31940
rect 3080 -32020 3100 -31960
rect 3160 -32020 3180 -31960
rect 3080 -32040 3180 -32020
rect 3880 -31960 3980 -31940
rect 3880 -32020 3900 -31960
rect 3960 -32020 3980 -31960
rect 3880 -32040 3980 -32020
rect 5480 -31960 5580 -31940
rect 5480 -32020 5500 -31960
rect 5560 -32020 5580 -31960
rect 5480 -32040 5580 -32020
rect -6260 -32104 -6220 -32040
rect -5460 -32104 -5420 -32040
rect -4660 -32104 -4620 -32040
rect -6268 -32148 -6212 -32104
rect -5468 -32148 -5412 -32104
rect -4668 -32148 -4612 -32104
rect -3860 -32120 -3820 -32040
rect -2260 -32100 -2220 -32040
rect -1460 -32100 -1420 -32040
rect 740 -32100 780 -32040
rect 1540 -32088 1580 -32040
rect 2340 -32088 2380 -32040
rect 3140 -32088 3180 -32040
rect 3940 -32088 3980 -32040
rect -2268 -32144 -2212 -32100
rect 1532 -32132 1588 -32088
rect 2332 -32132 2388 -32088
rect 3132 -32132 3188 -32088
rect 3932 -32132 3988 -32088
rect -6268 -32976 -6212 -32932
rect -5468 -32976 -5412 -32932
rect -4668 -32976 -4612 -32932
rect 5540 -32140 5580 -32040
rect 1532 -32736 1588 -32692
rect 2332 -32736 2388 -32692
rect 3132 -32736 3188 -32692
rect 3932 -32736 3988 -32692
rect -2268 -33720 -2212 -33712
rect -2268 -33756 -2260 -33720
rect -6344 -34173 -6144 -34160
rect -6344 -34219 -6331 -34173
rect -6157 -34219 -6144 -34173
rect -6344 -34282 -6144 -34219
rect -6344 -62345 -6144 -62282
rect -6344 -62391 -6331 -62345
rect -6157 -62391 -6144 -62345
rect -6344 -62404 -6144 -62391
rect -5544 -34173 -5344 -34160
rect -5544 -34219 -5531 -34173
rect -5357 -34219 -5344 -34173
rect -5544 -34282 -5344 -34219
rect -5544 -62345 -5344 -62282
rect -5544 -62391 -5531 -62345
rect -5357 -62391 -5344 -62345
rect -5544 -62404 -5344 -62391
rect -4744 -34173 -4544 -34160
rect -4744 -34219 -4731 -34173
rect -4557 -34219 -4544 -34173
rect -4744 -34282 -4544 -34219
rect -4744 -62345 -4544 -62282
rect -4744 -62391 -4731 -62345
rect -4557 -62391 -4544 -62345
rect -4744 -62404 -4544 -62391
rect -3944 -34173 -3744 -34160
rect -3944 -34219 -3931 -34173
rect -3757 -34219 -3744 -34173
rect -3944 -34282 -3744 -34219
rect -3944 -62345 -3744 -62282
rect -3944 -62391 -3931 -62345
rect -3757 -62391 -3744 -62345
rect -3944 -62404 -3744 -62391
rect -2344 -34180 -2260 -34160
rect -2160 -34180 -2144 -34160
rect -2344 -34282 -2144 -34180
rect -2344 -62345 -2144 -62282
rect -2344 -62391 -2331 -62345
rect -2157 -62391 -2144 -62345
rect -2344 -62404 -2144 -62391
rect -1544 -34173 -1344 -34160
rect -1544 -34219 -1531 -34173
rect -1357 -34219 -1344 -34173
rect -1544 -34282 -1344 -34219
rect -1544 -62345 -1344 -62282
rect -1544 -62391 -1531 -62345
rect -1357 -62391 -1344 -62345
rect -1544 -62404 -1344 -62391
rect 656 -34133 856 -34120
rect 656 -34179 669 -34133
rect 843 -34179 856 -34133
rect 656 -34242 856 -34179
rect 656 -62305 856 -62242
rect 656 -62351 669 -62305
rect 843 -62351 856 -62305
rect 656 -62364 856 -62351
rect 1456 -34133 1656 -34120
rect 1456 -34179 1469 -34133
rect 1643 -34179 1656 -34133
rect 1456 -34242 1656 -34179
rect 1456 -62305 1656 -62242
rect 1456 -62351 1469 -62305
rect 1643 -62351 1656 -62305
rect 1456 -62364 1656 -62351
rect 2256 -34133 2456 -34120
rect 2256 -34179 2269 -34133
rect 2443 -34179 2456 -34133
rect 2256 -34242 2456 -34179
rect 2256 -62305 2456 -62242
rect 2256 -62351 2269 -62305
rect 2443 -62351 2456 -62305
rect 2256 -62364 2456 -62351
rect 3056 -34133 3256 -34120
rect 3056 -34179 3069 -34133
rect 3243 -34179 3256 -34133
rect 3056 -34242 3256 -34179
rect 3056 -62305 3256 -62242
rect 3056 -62351 3069 -62305
rect 3243 -62351 3256 -62305
rect 3056 -62364 3256 -62351
rect 3856 -34133 4056 -34120
rect 3856 -34179 3869 -34133
rect 4043 -34179 4056 -34133
rect 3856 -34242 4056 -34179
rect 3856 -62305 4056 -62242
rect 3856 -62351 3869 -62305
rect 4043 -62351 4056 -62305
rect 3856 -62364 4056 -62351
rect 5456 -34133 5656 -34120
rect 5456 -34179 5469 -34133
rect 5643 -34179 5656 -34133
rect 5456 -34242 5656 -34179
rect 5456 -62305 5656 -62242
rect 5456 -62351 5469 -62305
rect 5643 -62351 5656 -62305
rect 5456 -62364 5656 -62351
<< polycontact >>
rect -5580 -820 -5500 -740
rect -520 -820 -440 -740
rect -160 -820 -80 -740
rect 4900 -820 4980 -740
rect -5580 -1260 -5500 -1180
rect 4916 -1260 4996 -1180
rect -9940 -2060 -9880 -2000
rect -9600 -2060 -9540 -2000
rect 6180 -2820 6240 -2760
rect 6180 -2980 6240 -2920
rect -6331 -3519 -6157 -3473
rect -6331 -31691 -6157 -31645
rect -5531 -3519 -5357 -3473
rect -5531 -31691 -5357 -31645
rect -4731 -3519 -4557 -3473
rect -4731 -31691 -4557 -31645
rect -3931 -3519 -3757 -3473
rect -3931 -31691 -3757 -31645
rect -2331 -3519 -2157 -3473
rect -2331 -31691 -2157 -31645
rect -1531 -3519 -1357 -3473
rect -1531 -31691 -1357 -31645
rect 1469 -3519 1643 -3473
rect 1469 -31691 1643 -31645
rect 2269 -3519 2443 -3473
rect 2269 -31691 2443 -31645
rect 3069 -3519 3243 -3473
rect 3069 -31691 3243 -31645
rect 3869 -3519 4043 -3473
rect 3869 -31691 4043 -31645
rect 5469 -3519 5643 -3473
rect 5469 -31691 5643 -31645
rect -6240 -32020 -6180 -31960
rect -5440 -32020 -5380 -31960
rect -4640 -32020 -4580 -31960
rect -3840 -32020 -3780 -31960
rect -2240 -32020 -2180 -31960
rect -1440 -32020 -1380 -31960
rect 700 -32020 760 -31960
rect 1500 -32020 1560 -31960
rect 2300 -32020 2360 -31960
rect 3100 -32020 3160 -31960
rect 3900 -32020 3960 -31960
rect 5500 -32020 5560 -31960
rect -6331 -34219 -6157 -34173
rect -6331 -62391 -6157 -62345
rect -5531 -34219 -5357 -34173
rect -5531 -62391 -5357 -62345
rect -4731 -34219 -4557 -34173
rect -4731 -62391 -4557 -62345
rect -3931 -34219 -3757 -34173
rect -3931 -62391 -3757 -62345
rect -2331 -62391 -2157 -62345
rect -1531 -34219 -1357 -34173
rect -1531 -62391 -1357 -62345
rect 669 -34179 843 -34133
rect 669 -62351 843 -62305
rect 1469 -34179 1643 -34133
rect 1469 -62351 1643 -62305
rect 2269 -34179 2443 -34133
rect 2269 -62351 2443 -62305
rect 3069 -34179 3243 -34133
rect 3069 -62351 3243 -62305
rect 3869 -34179 4043 -34133
rect 3869 -62351 4043 -62305
rect 5469 -34179 5643 -34133
rect 5469 -62351 5643 -62305
<< nhighres >>
rect -6344 -31582 -6144 -3582
rect -5544 -31582 -5344 -3582
rect -4744 -31582 -4544 -3582
rect -3944 -31582 -3744 -3582
rect -2344 -31582 -2144 -3582
rect -1544 -31582 -1344 -3582
rect 1456 -31582 1656 -3582
rect 2256 -31582 2456 -3582
rect 3056 -31582 3256 -3582
rect 3856 -31582 4056 -3582
rect 5456 -31582 5656 -3582
rect -6344 -62282 -6144 -34282
rect -5544 -62282 -5344 -34282
rect -4744 -62282 -4544 -34282
rect -3944 -62282 -3744 -34282
rect -2344 -62282 -2144 -34282
rect -1544 -62282 -1344 -34282
rect 656 -62242 856 -34242
rect 1456 -62242 1656 -34242
rect 2256 -62242 2456 -34242
rect 3056 -62242 3256 -34242
rect 3856 -62242 4056 -34242
rect 5456 -62242 5656 -34242
<< pdiffres >>
rect -1768 66 -848 266
<< metal1 >>
rect -1881 253 -1835 264
rect -3220 80 -1881 240
rect -3220 -380 -3140 80
rect -380 240 -220 760
rect -780 80 180 240
rect 1280 80 2640 240
rect -1881 68 -1835 79
rect -5780 -400 -3140 -380
rect 2560 -220 2640 80
rect 2620 -300 2640 -220
rect -5780 -480 140 -400
rect -5780 -500 -3140 -480
rect -3220 -680 -3140 -500
rect -760 -560 -640 -540
rect -760 -620 -740 -560
rect -660 -620 -640 -560
rect -760 -680 -640 -620
rect -720 -720 -640 -680
rect -360 -560 -240 -540
rect -360 -620 -340 -560
rect -260 -620 -240 -560
rect -360 -740 -240 -620
rect 60 -677 140 -480
rect 2560 -677 2640 -300
rect 50 -723 61 -677
rect 2275 -723 2286 -677
rect 2550 -723 2561 -677
rect 4775 -723 4786 -677
rect -5780 -820 -5580 -740
rect -5500 -820 -5480 -740
rect -540 -820 -520 -740
rect -440 -820 -160 -740
rect -80 -820 -60 -740
rect 4880 -820 4900 -740
rect 4980 -820 5180 -740
rect -5360 -1160 -5280 -840
rect -980 -1160 -900 -840
rect 50 -883 61 -837
rect 2275 -883 2286 -837
rect 2550 -883 2561 -837
rect 4775 -883 4786 -837
rect 320 -1120 400 -883
rect 4700 -1120 4780 -883
rect -5780 -1260 -5580 -1180
rect -5500 -1260 -5480 -1180
rect 4896 -1260 4916 -1180
rect 4996 -1260 5196 -1180
rect -940 -1340 -880 -1280
rect 300 -1340 360 -1280
rect -940 -1400 360 -1340
rect -14100 -1860 -9700 -1780
rect -14100 -2180 -13920 -1860
rect -13400 -1957 -10060 -1860
rect -13410 -2003 -13399 -1957
rect -10065 -2003 -10054 -1957
rect -9780 -1980 -9700 -1860
rect -6140 -1880 -2960 -1800
rect -6140 -1960 -6060 -1880
rect -9960 -2000 -9520 -1980
rect -9960 -2060 -9940 -2000
rect -9880 -2060 -9600 -2000
rect -9540 -2060 -9520 -2000
rect -9960 -2080 -9520 -2060
rect -13410 -2163 -13399 -2117
rect -10065 -2140 -10054 -2117
rect -10065 -2163 -9360 -2140
rect -10100 -2200 -9360 -2163
rect -5080 -2940 -5000 -2920
rect -5080 -3000 -5060 -2940
rect -5080 -3460 -5000 -3000
rect -6340 -3473 -3740 -3460
rect -6342 -3519 -6331 -3473
rect -6157 -3519 -5531 -3473
rect -5357 -3519 -4731 -3473
rect -4557 -3519 -3931 -3473
rect -3757 -3519 -3740 -3473
rect -6340 -3520 -3740 -3519
rect -14100 -3920 -7020 -3840
rect -7180 -32160 -7020 -3920
rect -6260 -31645 -6160 -31640
rect -5460 -31645 -5360 -31640
rect -4660 -31645 -4560 -31640
rect -3860 -31645 -3760 -31640
rect -6342 -31691 -6331 -31645
rect -6157 -31691 -6146 -31645
rect -5542 -31691 -5531 -31645
rect -5357 -31691 -5346 -31645
rect -4742 -31691 -4731 -31645
rect -4557 -31691 -4546 -31645
rect -3942 -31691 -3931 -31645
rect -3757 -31691 -3746 -31645
rect -6260 -31960 -6160 -31691
rect -6260 -32020 -6240 -31960
rect -6180 -32020 -6160 -31960
rect -6260 -32040 -6160 -32020
rect -5460 -31960 -5360 -31691
rect -5460 -32020 -5440 -31960
rect -5380 -32020 -5360 -31960
rect -5460 -32040 -5360 -32020
rect -4660 -31960 -4560 -31691
rect -4660 -32020 -4640 -31960
rect -4580 -32020 -4560 -31960
rect -4660 -32040 -4560 -32020
rect -3860 -31960 -3760 -31691
rect -3860 -32020 -3840 -31960
rect -3780 -32020 -3760 -31960
rect -3860 -32040 -3760 -32020
rect -6343 -32160 -6297 -32150
rect -7180 -32161 -6297 -32160
rect -7180 -32320 -6343 -32161
rect -7180 -34480 -7020 -32320
rect -6343 -32930 -6297 -32919
rect -6183 -32160 -6137 -32150
rect -5543 -32160 -5497 -32150
rect -6183 -32161 -5497 -32160
rect -6137 -32919 -5543 -32161
rect -6183 -32920 -5497 -32919
rect -6183 -32930 -6137 -32920
rect -5543 -32930 -5497 -32920
rect -5383 -32160 -5337 -32150
rect -4743 -32160 -4697 -32150
rect -5383 -32161 -4697 -32160
rect -5337 -32919 -4743 -32161
rect -5383 -32920 -4697 -32919
rect -5383 -32930 -5337 -32920
rect -4743 -32930 -4697 -32920
rect -4583 -32160 -4537 -32150
rect -3120 -32160 -2960 -1880
rect -1880 -3120 -1800 -3100
rect -1880 -3180 -1860 -3120
rect -1880 -3460 -1800 -3180
rect -2340 -3473 -1340 -3460
rect -2342 -3519 -2331 -3473
rect -2157 -3519 -1531 -3473
rect -1357 -3519 -1340 -3473
rect -2340 -3520 -1340 -3519
rect -2260 -31645 -2160 -31640
rect -1460 -31645 -1360 -31640
rect -2342 -31691 -2331 -31645
rect -2157 -31691 -2146 -31645
rect -1542 -31691 -1531 -31645
rect -1357 -31691 -1346 -31645
rect -2260 -31960 -2160 -31691
rect -2260 -32020 -2240 -31960
rect -2180 -32020 -2160 -31960
rect -2260 -32040 -2160 -32020
rect -1460 -31960 -1360 -31691
rect -1460 -32020 -1440 -31960
rect -1380 -32020 -1360 -31960
rect -1460 -32040 -1360 -32020
rect -380 -32140 -220 -1400
rect 4700 -1940 6860 -1780
rect 2320 -2940 2400 -2920
rect 2380 -3000 2400 -2940
rect 2320 -3460 2400 -3000
rect 660 -3473 4060 -3460
rect 660 -3519 1469 -3473
rect 1643 -3519 2269 -3473
rect 2443 -3519 3069 -3473
rect 3243 -3519 3869 -3473
rect 4043 -3519 4060 -3473
rect 660 -3520 4060 -3519
rect 680 -31960 780 -31640
rect 1480 -31645 1580 -31640
rect 2280 -31645 2380 -31640
rect 3080 -31645 3180 -31640
rect 3880 -31645 3980 -31640
rect 1458 -31691 1469 -31645
rect 1643 -31691 1654 -31645
rect 2258 -31691 2269 -31645
rect 2443 -31691 2454 -31645
rect 3058 -31691 3069 -31645
rect 3243 -31691 3254 -31645
rect 3858 -31691 3869 -31645
rect 4043 -31691 4054 -31645
rect 680 -32020 700 -31960
rect 760 -32020 780 -31960
rect 680 -32040 780 -32020
rect 1480 -31960 1580 -31691
rect 1480 -32020 1500 -31960
rect 1560 -32020 1580 -31960
rect 1480 -32040 1580 -32020
rect 2280 -31960 2380 -31691
rect 2280 -32020 2300 -31960
rect 2360 -32020 2380 -31960
rect 2280 -32040 2380 -32020
rect 3080 -31960 3180 -31691
rect 3080 -32020 3100 -31960
rect 3160 -32020 3180 -31960
rect 3080 -32040 3180 -32020
rect 3880 -31960 3980 -31691
rect 3880 -32020 3900 -31960
rect 3960 -32020 3980 -31960
rect 3880 -32040 3980 -32020
rect 1457 -32140 1503 -32134
rect -2343 -32157 -2297 -32146
rect -4583 -32161 -3900 -32160
rect -4537 -32919 -3900 -32161
rect -4583 -32920 -3900 -32919
rect -3780 -32920 -2343 -32160
rect -4583 -32930 -4537 -32920
rect -2343 -33710 -2297 -33699
rect -2183 -32157 -2137 -32146
rect -2137 -33699 -1500 -32160
rect -1340 -32680 700 -32140
rect 820 -32145 1503 -32140
rect 820 -32679 1457 -32145
rect 820 -32680 1503 -32679
rect 1457 -32690 1503 -32680
rect 1617 -32140 1663 -32134
rect 2257 -32140 2303 -32134
rect 1617 -32145 2303 -32140
rect 1663 -32679 2257 -32145
rect 1617 -32680 2303 -32679
rect 1617 -32690 1663 -32680
rect 2257 -32690 2303 -32680
rect 2417 -32140 2463 -32134
rect 3057 -32140 3103 -32134
rect 2417 -32145 3103 -32140
rect 2463 -32679 3057 -32145
rect 2417 -32680 3103 -32679
rect 2417 -32690 2463 -32680
rect 3057 -32690 3103 -32680
rect 3217 -32140 3263 -32134
rect 3857 -32140 3903 -32134
rect 3217 -32145 3903 -32140
rect 3263 -32679 3857 -32145
rect 3217 -32680 3903 -32679
rect 3217 -32690 3263 -32680
rect 3857 -32690 3903 -32680
rect 4017 -32140 4063 -32134
rect 4700 -32140 4860 -1940
rect 6100 -2220 6200 -2200
rect 6100 -2280 6120 -2220
rect 6180 -2280 6200 -2220
rect 6100 -2300 6200 -2280
rect 6120 -2600 6180 -2300
rect 6300 -2640 6360 -2440
rect 6300 -2680 6380 -2640
rect 6160 -2760 6260 -2740
rect 6160 -2820 6180 -2760
rect 6240 -2820 6260 -2760
rect 5500 -2840 5600 -2820
rect 6160 -2840 6260 -2820
rect 5500 -2900 5520 -2840
rect 5580 -2900 6260 -2840
rect 5500 -2920 5600 -2900
rect 6160 -2920 6260 -2900
rect 6160 -2980 6180 -2920
rect 6240 -2980 6260 -2920
rect 6160 -3000 6260 -2980
rect 6320 -2820 6380 -2680
rect 6320 -2840 6520 -2820
rect 6320 -2900 6440 -2840
rect 6500 -2900 6520 -2840
rect 6320 -2920 6520 -2900
rect 6320 -3080 6380 -2920
rect 5520 -3120 5600 -3100
rect 5580 -3180 5600 -3120
rect 5520 -3473 5600 -3180
rect 5458 -3519 5469 -3473
rect 5643 -3519 5654 -3473
rect 5520 -3520 5600 -3519
rect 6120 -3620 6180 -3100
rect 6300 -3120 6380 -3080
rect 6300 -3260 6360 -3120
rect 5480 -31645 5580 -31640
rect 5458 -31691 5469 -31645
rect 5643 -31691 5654 -31645
rect 5480 -31960 5580 -31691
rect 5480 -32020 5500 -31960
rect 5560 -32020 5580 -31960
rect 5480 -32040 5580 -32020
rect 4017 -32145 5500 -32140
rect 4063 -32300 5500 -32145
rect 5620 -32300 6340 -32140
rect 4017 -32690 4063 -32679
rect -2183 -33700 -1500 -33699
rect 6180 -33340 6340 -32300
rect 6180 -33500 6940 -33340
rect -2183 -33710 -2137 -33700
rect -6280 -34160 -6200 -33820
rect -5480 -34160 -5400 -33820
rect -4680 -34160 -4600 -33820
rect -3880 -34160 -3800 -33820
rect -6280 -34173 -6160 -34160
rect -5480 -34173 -5360 -34160
rect -4680 -34173 -4560 -34160
rect -3880 -34173 -3760 -34160
rect -6342 -34219 -6331 -34173
rect -6157 -34219 -6146 -34173
rect -5542 -34219 -5531 -34173
rect -5357 -34219 -5346 -34173
rect -4742 -34219 -4731 -34173
rect -4557 -34219 -4546 -34173
rect -3942 -34219 -3931 -34173
rect -3757 -34219 -3746 -34173
rect -2280 -34180 -2200 -33760
rect -1480 -34160 -1400 -33760
rect 720 -34120 800 -33780
rect 1520 -34120 1600 -33780
rect 2320 -34120 2400 -33780
rect 3120 -34120 3200 -33780
rect 3920 -34120 4000 -33780
rect 5520 -34120 5600 -33780
rect 720 -34133 840 -34120
rect 1520 -34133 1640 -34120
rect 2320 -34133 2440 -34120
rect 3120 -34133 3240 -34120
rect 3920 -34133 4040 -34120
rect 5520 -34133 5640 -34120
rect -1480 -34173 -1360 -34160
rect -6260 -34220 -6160 -34219
rect -5460 -34220 -5360 -34219
rect -4660 -34220 -4560 -34219
rect -3860 -34220 -3760 -34219
rect -2260 -34220 -2160 -34180
rect -1542 -34219 -1531 -34173
rect -1357 -34219 -1346 -34173
rect 658 -34179 669 -34133
rect 843 -34179 854 -34133
rect 1458 -34179 1469 -34133
rect 1643 -34179 1654 -34133
rect 2258 -34179 2269 -34133
rect 2443 -34179 2454 -34133
rect 3058 -34179 3069 -34133
rect 3243 -34179 3254 -34133
rect 3858 -34179 3869 -34133
rect 4043 -34179 4054 -34133
rect 5458 -34179 5469 -34133
rect 5643 -34179 5654 -34133
rect 740 -34180 840 -34179
rect 1540 -34180 1640 -34179
rect 2340 -34180 2440 -34179
rect 3140 -34180 3240 -34179
rect 3940 -34180 4040 -34179
rect 5540 -34180 5640 -34179
rect -1460 -34220 -1360 -34219
rect 6180 -34480 6340 -33500
rect -7180 -34640 6340 -34480
rect 740 -62305 840 -62300
rect 1540 -62305 1640 -62300
rect 2340 -62305 2440 -62300
rect 3140 -62305 3240 -62300
rect 3940 -62305 4040 -62300
rect 5540 -62305 5640 -62300
rect -6260 -62345 -6160 -62340
rect -5460 -62345 -5360 -62340
rect -4660 -62345 -4560 -62340
rect -3860 -62345 -3760 -62340
rect -2260 -62345 -2160 -62340
rect -1460 -62345 -1360 -62340
rect -6342 -62391 -6331 -62345
rect -6157 -62391 -6146 -62345
rect -5542 -62391 -5531 -62345
rect -5357 -62391 -5346 -62345
rect -4742 -62391 -4731 -62345
rect -4557 -62391 -4546 -62345
rect -3942 -62391 -3931 -62345
rect -3757 -62391 -3746 -62345
rect -2342 -62391 -2331 -62345
rect -2157 -62391 -2146 -62345
rect -1542 -62391 -1531 -62345
rect -1357 -62391 -1346 -62345
rect 658 -62351 669 -62305
rect 843 -62351 854 -62305
rect 1458 -62351 1469 -62305
rect 1643 -62351 1654 -62305
rect 2258 -62351 2269 -62305
rect 2443 -62351 2454 -62305
rect 3058 -62351 3069 -62305
rect 3243 -62351 3254 -62305
rect 3858 -62351 3869 -62305
rect 4043 -62351 4054 -62305
rect 5458 -62351 5469 -62305
rect 5643 -62351 5654 -62305
rect -6260 -62680 -6160 -62391
rect -5460 -62680 -5360 -62391
rect -4660 -62680 -4560 -62391
rect -3860 -62680 -3760 -62391
rect -2260 -62680 -2160 -62391
rect -1460 -62680 -1360 -62391
rect 740 -62680 840 -62351
rect 1540 -62680 1640 -62351
rect 2340 -62680 2440 -62351
rect 3140 -62680 3240 -62351
rect 3940 -62680 4040 -62351
rect 5540 -62680 5640 -62351
rect -6560 -62840 6660 -62680
<< via1 >>
rect 2560 -300 2620 -220
rect -740 -620 -660 -560
rect -340 -620 -260 -560
rect -5060 -3000 -5000 -2940
rect -1860 -3180 -1800 -3120
rect 2320 -3000 2380 -2940
rect 6120 -2280 6180 -2220
rect 5520 -2900 5580 -2840
rect 6440 -2900 6500 -2840
rect 5520 -3180 5580 -3120
<< metal2 >>
rect -760 -220 5180 -200
rect -760 -300 2560 -220
rect 2620 -300 5180 -220
rect -760 -320 5180 -300
rect -760 -560 -640 -320
rect -760 -620 -740 -560
rect -660 -620 -640 -560
rect -760 -640 -640 -620
rect -360 -560 5180 -540
rect -360 -620 -340 -560
rect -260 -620 5180 -560
rect -360 -640 5180 -620
rect 5500 -2140 6860 -2040
rect 5500 -2840 5600 -2140
rect 6100 -2220 6860 -2200
rect 6100 -2280 6120 -2220
rect 6180 -2280 6860 -2220
rect 6100 -2300 6860 -2280
rect 5500 -2900 5520 -2840
rect 5580 -2900 5600 -2840
rect 5500 -2920 5600 -2900
rect -5080 -2940 5600 -2920
rect -5080 -3000 -5060 -2940
rect -5000 -3000 2320 -2940
rect 2380 -3000 5600 -2940
rect -5080 -3020 5600 -3000
rect 6420 -2840 6520 -2820
rect 6420 -2900 6440 -2840
rect 6500 -2900 6520 -2840
rect -1880 -3120 6020 -3100
rect -1880 -3180 -1860 -3120
rect -1800 -3180 5520 -3120
rect 5580 -3180 6020 -3120
rect -1880 -3200 6020 -3180
rect 5920 -3420 6020 -3200
rect 6420 -3420 6520 -2900
rect 5920 -3520 6520 -3420
use nfet_03v3_EF5H4U  nfet_03v3_EF5H4U_0
timestamp 1757524825
transform 1 0 6240 0 1 -3184
box -140 -156 140 156
use nfet_03v3_N5W335  nfet_03v3_N5W335_0
timestamp 1757529591
transform 1 0 -1440 0 1 -32928
box -140 -852 140 852
use nfet_03v3_N5W335  nfet_03v3_N5W335_1
timestamp 1757529591
transform 1 0 -2240 0 1 -32928
box -140 -852 140 852
use nfet_03v3_N5WHL5  nfet_03v3_N5WHL5_0
timestamp 1757529591
transform 1 0 5560 0 1 -32228
box -140 -152 140 152
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_0
timestamp 1757529591
transform 1 0 -3840 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_1
timestamp 1757529591
transform 1 0 -4640 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_2
timestamp 1757529591
transform 1 0 -6240 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NL3C35  nfet_03v3_NL3C35_3
timestamp 1757529591
transform 1 0 -5440 0 1 -32540
box -140 -460 140 460
use nfet_03v3_NMLPX4  nfet_03v3_NMLPX4_0
timestamp 1757063525
transform 0 1 -3132 -1 0 -1220
box -140 -2308 140 2308
use nfet_03v3_NMLPX4  nfet_03v3_NMLPX4_1
timestamp 1757063525
transform 0 1 2548 -1 0 -1220
box -140 -2308 140 2308
use nfet_03v3_NP3335  nfet_03v3_NP3335_0
timestamp 1757535309
transform 0 1 -7732 -1 0 -2060
box -140 -1748 140 1748
use nfet_03v3_NP3335  nfet_03v3_NP3335_1
timestamp 1757535309
transform 0 1 -11732 -1 0 -2060
box -140 -1748 140 1748
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_0
timestamp 1757527981
transform 1 0 760 0 1 -32412
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_1
timestamp 1757527981
transform 1 0 1560 0 1 -32412
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_2
timestamp 1757527981
transform 1 0 2360 0 1 -32412
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_3
timestamp 1757527981
transform 1 0 3160 0 1 -32412
box -140 -348 140 348
use nfet_03v3_NPKKZ4  nfet_03v3_NPKKZ4_4
timestamp 1757527981
transform 1 0 3960 0 1 -32412
box -140 -348 140 348
use nfet_03v3_NUG935  nfet_03v3_NUG935_0
timestamp 1757012598
transform 0 1 -4252 -1 0 -780
box -140 -1188 140 1188
use nfet_03v3_NUG935  nfet_03v3_NUG935_1
timestamp 1757012598
transform 0 1 -1752 -1 0 -780
box -140 -1188 140 1188
use nfet_03v3_NUG935  nfet_03v3_NUG935_2
timestamp 1757012598
transform 0 1 3668 -1 0 -780
box -140 -1188 140 1188
use nfet_03v3_NUG935  nfet_03v3_NUG935_3
timestamp 1757012598
transform 0 1 1168 -1 0 -780
box -140 -1188 140 1188
use pfet_03v3_6ZJ338  pfet_03v3_6ZJ338_0
timestamp 1757524825
transform 1 0 6242 0 1 -2522
box -202 -218 202 218
use pplus_u_CRD77H  pplus_u_CRD77H_0
timestamp 1757010180
transform 0 1 712 -1 0 166
box -286 -772 286 772
use pplus_u_CRD77H  pplus_u_CRD77H_1
timestamp 1757010180
transform 0 -1 -1308 1 0 166
box -286 -772 286 772
use ppolyf_u_1k_4GNJYW  ppolyf_u_1k_4GNJYW_0
timestamp 1757535624
transform 1 0 -14004 0 1 -3032
box -336 -1108 336 1108
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_0
timestamp 1757065516
transform 1 0 756 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_1
timestamp 1757065516
transform 1 0 1556 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_2
timestamp 1757065516
transform 1 0 2356 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_3
timestamp 1757065516
transform 1 0 3156 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_4
timestamp 1757065516
transform 1 0 3956 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_5
timestamp 1757065516
transform 1 0 5556 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_6
timestamp 1757065516
transform 1 0 -1444 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_7
timestamp 1757065516
transform 1 0 -2244 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_8
timestamp 1757065516
transform 1 0 -3844 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_9
timestamp 1757065516
transform 1 0 -5444 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_10
timestamp 1757065516
transform 1 0 -6244 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_11
timestamp 1757065516
transform 1 0 -4644 0 1 -17582
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_12
timestamp 1757065516
transform 1 0 -2244 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_13
timestamp 1757065516
transform 1 0 -1444 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_14
timestamp 1757065516
transform 1 0 756 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_15
timestamp 1757065516
transform 1 0 1556 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_16
timestamp 1757065516
transform 1 0 2356 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_17
timestamp 1757065516
transform 1 0 3156 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_18
timestamp 1757065516
transform 1 0 3956 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_19
timestamp 1757065516
transform 1 0 5556 0 1 -48242
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_20
timestamp 1757065516
transform 1 0 -3844 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_21
timestamp 1757065516
transform 1 0 -4644 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_22
timestamp 1757065516
transform 1 0 -5444 0 1 -48282
box -336 -14358 336 14358
use ppolyf_u_1k_9FJPHG  ppolyf_u_1k_9FJPHG_23
timestamp 1757065516
transform 1 0 -6244 0 1 -48282
box -336 -14358 336 14358
<< end >>
